library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;



entity table_3000 is


    Port ( Clk   : in std_logic;
           ADDR  : in integer  range 0 to 1023; 
           DOUT  : out integer range 0 to 999999;
           LOUT  : out integer range 0 to 1 
	);

end table_3000;

architecture Behavioral of table_3000 is
type matrice_angulo3000 is array (0 to 115) of integer range 0 to 999999;  
type matrice_bit3000    is array (0 to 115) of integer range 0 to 1; 

constant angulos3000: matrice_angulo3000 :=( 

-- ************ Ma=0.8 ************* --
15998 	,
17394 	,
32002 	,
34779 	,
48019 	,
52146 	,
64056 	,
69486 	,
80118 	,
86792 	,
96211 	,
104055	,
112342	,
121269	,
128517	,
138428	,
144739	,
155527	,
161015	,
172560	,
177350	,
189525	,
193746	,
206419	,
210208	,
223240	,
226738	,
239987	,
243339	,
256661	,
260013	,
273262	,
276760	,
289792	,
293581	,
306254	,
310475	,
322650	,
327440	,
338985	,
344473	,
355261	,
361572	,
371483	,
378731	,
387658	,
395945	,
403789	,
413208	,
419882	,
430514	,
435944	,
447854	,
451981	,
465221	,
467998	,
482606	,
484002	,
515998	,
517394	,
532002	,
534779	,
548019	,
552146	,
564056	,
569486	,
580118	,
586792	,
596211	,
604055	,
612342	,
621269	,
628517	,
638428	,
644739	,
655527	,
661015	,
672560	,
677350	,
689525	,
693746	,
706419	,
710208	,
723240	,
726738	,
739987	,
743339	,
756661	,
760013	,
773262	,
776760	,
789792	,
793581	,
806254	,
810475	,
822650	,
827440	,
838985	,
844473	,
855261	,
861572	,
871483	,
878731	,
887658	,
895945	,
903789	,
913208	,
919882	,
930514	,
935944	,
947854	,
951981	,
965221	,
967998	,
982606	,
984002	
      	
	
      



            
-- ******************************** --
);

constant nivel3000: matrice_bit3000 :=( 

-- ************ Ma=0.8 ************* --
0       ,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	,
0	,
1	




	


            
-- ******************************** --
);


begin
  Process(Clk)
    begin 
      if Clk'event and Clk='1' then
         DOUT <= angulos3000(ADDR);
         LOUT <= nivel3000(ADDR);
      end if;
  end process;
      
end Behavioral;



